/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	oops_assign3.sv  
Date:   	30th May 2024
Version:	1.0
Description: Concept of OOPS in SV 
***************************************************************************/
class base;
  //ADD_CODE: Add a void vitrual function with the name display();
  //ADD_CODE: Display a string with the name of the base class $display ("base_class);
endclass

//ADD_CODE: Extend the base class with a name derived class 
  //ADD_CODE: To overide the method of the base class 
  //ADD_CODE: Add the function with the same name mentioned in the base class and use the OOPS principle to override 
  //ADD_CODE: Display the string with the name of the derived class 
endclass

module poly;
initial  
  begin
    //ADD_CODE: To create the instances and object of base class
    //ADD_CODE: To create the instances and object of derived class

    //ADD_CODE: Call the display method of the base class 
    //ADD_CODE: Call the display method of derived class 

    //ADD_CODE: Do a simple copy to point the instance of base class to derived class object
    //ADD_CODE: Call the display method of the base class 
    //ADD_CODE: Call the display method of derived class 
  end
endmodule



