/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	func_assign1.sv  
Date:   	7th June 2024
Version:	1.0
Description: Concept of Caonstraint Randomization in System Verilog 
***************************************************************************/
class constraint_assign1;
  
//ADD_CODE: Declare the 8bit variable as data. 
//ADD_CODE: Write constraint for an 8bit variable data to generate values divisible by 5.
  
endclass
module con_assin1; 
initial
  begin
    //ADD_CODE: Call the function addition and pass the argument by value
    //Return the value of the function  by using a return statement 
    //ADD_CODE: Display the values of the result
    
    //ADD_CODE: Call the function addition and pass the argument by 
    //Return the value by assigning a value to the internal variable with the same name as the function
    //ADD_CODE: Display the values of the result
    

  end
endmodule
