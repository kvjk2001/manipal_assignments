/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	data_assign4.sv  
Date:   	21st May 2022
Version:	1.0
Description: Concept of structure data type 
***************************************************************************/
//Declare the struct with name money as typedef
//Store coins as type int and rupees as real

module data_assign4;
 //To create the instance of the structure
  initial 
    begin
      //Assign directvalues to the structure variables
      //Display the values of the memebers
    
      //Assign values using the memebers name
      //Display the values 
    
      //Assign all elements of structure to zero
      //Display the values 
  end
endmodule
