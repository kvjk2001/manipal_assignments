/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	data_assign2.sv  
Date:   	21st May 2022
Version:	1.0
Description: Concept of associative array and functions 
***************************************************************************/
// Write a function to return a dynamic array of size 10 filled with random integers.
module data_assign2;

  //Part 1
  //ADD_CODE: Declare a function and input the size 
  //ADD_CODE: Inside the function declare and create the array
  //ADD_CODE: Use the appropriate loop to randomize the elemants of the array


  //Part 2a
  //ADD_CODE: The array method to return the maximum value stored in the array


  //part 2b
  //ADD_CODE: Modify the Part 1 function to arrange the array with out array method
  //ADD_CODE: write a function to arrange the the array in the ascending order
  //HINT : using a loop you can compare the values of the array with previous value
  

  initial 
    begin
      repeat(30)
      //ADD_CODE: call the function
      //ADD_CODE: Display the elements of the dynamic array
      //ADD_CODE: Display the array and the maximum value 
      //ADD_CODE: Display the maximum value of the array and second largest value in the array
  
    end
endmodule
