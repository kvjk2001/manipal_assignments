/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	oops_assign5.sv  
Date:   	30th May 2024
Version:	1.0
Description: Write a code for an example of Shallow copy and Deep Copy 
***************************************************************************/
