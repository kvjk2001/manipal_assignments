/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	func_assign2.sv  
Date:   	7th June 2024
Version:	1.0
Description: Concept of Constraint Randomization in System Verilog 
***************************************************************************/
class constraint_assign2;
  
//ADD_CODE: Declare the 8bit variable as data. 
//ADD_CODE: Write constraint for a dynamic array address of size 10 to generate even numbers.
  
endclass:constraint_assign2 
module con_assin2; 
  //ADD_CODE: Declare the handle for "class constraint_assign2" as c0.
initial
  begin
    //ADD_CODE: Create the Object for  handle
    //ADD_CODE: Randomize the object for genrating randomize values for address with even numbers.
    //ADD_CODE: Display the values of of array address using object handel.
        
  end 
endmodule:con_assign2
