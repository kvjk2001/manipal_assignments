/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	data_assign2.sv  
Date:   	21st May 2022
Version:	1.0
Description: Concept of associative array and functions 
***************************************************************************/
// Write a function to return a dynamic array of size 10 filled with random integers.
module data_assign2;

  //Part 1
  //ADD_CODE: Declare a function and input the size 
  //ADD_CODE: Inside the function declare and create the array
  //ADD_CODE: Use the appropriate loop to randomize the elemants and display them

  //Part 2a
  //ADD_CODE: The array method to return the maximum value stored in the array
  //ADD_CODE: Display the array and the maximum value 

  //part 2b
  //ADD_CODE: Modify the Part 1 function to arrange the array with out array method
  //ADD_CODE: Display the maximum value of the array and the array 

  //Part 3
  //ADD_CODE: Display the second highest value 
  
  initial 
    begin
    repeat(30)
    //ADD_CODE: call the function
  end
endmodule
