/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	func_assign7.sv  
Date:   	7th June 2024
Version:	1.0
Description: Concept of Constraint Randomization in System Verilog 
***************************************************************************/
class constraint_assign7;
  
//ADD_CODE: Declare the 32bit variable. 
//ADD_CODE: Write for constraint to Generate a random 32-bit value With alternate pattern {0,1,0,1,...}  
  
endclass:constraint_assign7
module con_assin7; 
  //ADD_CODE: Declare the handle for "class constraint_assign7" as c0.
initial
  begin
    //ADD_CODE: Create the Object for  handle
          //ADD_CODE: Randomize the object for genrating randomize values of variable with pattern {0,1,0,1..}.
    //ADD_CODE: Display the values of variable using object handel.
        
  end 
endmodule:con_assign7
