/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	data_assign8.sv  
Date:   	21st May 2022
Version:	1.0
Description: Concept of associative array and dynamic array differences
***************************************************************************/
module data_assign8 (); // module name and file name same
  
  //ADD_CODE: Declare a dynamic array of dyn_arr
  //ADD_CODE: Declare the the size of an array
  //ADD_CODE: write a function to assign even values to the first 50 elements of the array
  //ADD_CODE: Display the value of the array 
  //ADD_CODE: Now write another function to add odd values to the last 50 elements 
  //ADD_CODE: Display all the 100 elements of the array
  //ADD_CODE: Write a method to delete the 90th element of the array
  //ADD_CODE: Write a method to delete the compelte array

  //Please repeat the same code with associative array with name assoc_arr and compare your findings
endmodule
 
