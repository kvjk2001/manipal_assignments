/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	func_assign9.sv  
Date:   	7th June 2024
Version:	1.0
Description: Concept of Constraint Randomization in System Verilog 
***************************************************************************/
class constraint_assign9;
  
//ADD_CODE: Declare the dynamic array fibo.
//ADD_CODE: Write for constraint to generate Fibonacci series.Ex: ( 0, 1, 1, 2, 3, 5, 8, 13, 21, 34, 55)

  
endclass:constraint_assign9
module con_assin9; 
  //ADD_CODE: Declare the handle for "class constraint_assign9" as c0.
initial
  begin
    //ADD_CODE: Create the Object for  handle
          //ADD_CODE: Randomize the object for genrating randomize values of array .
    //ADD_CODE: Display the values of array fibo  using object handel.
        
  end 
endmodule:con_assign9
