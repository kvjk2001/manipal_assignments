/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	oops_assign1.sv  
Date:   	22nd May 2024
Version:	1.0
Description: Concept of class constructor function and creation of Objects
***************************************************************************/
class construct
  //ADD_CODE: Declare a variable "i" of type int 
  //ADD_CODE: Decalre a class constructor function
endclass:construct

module class_cons;
  //ADD_CODE: declare the three handles c0,c1,c2 for the calss "construct"
initial
  begin
    //ADD_CODE: Create the Object for each handlle
    //ADD_CODE: Display the values of i for each object by using the class handle
    //ADD_CODE: Increment the value of "i" by 2  
    //ADD_CODE: Display the values of i for each object by using the class handle      
  end 
endmodule:class_cons
