/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	data_assign9.sv  
Date:   	24th May 2024
Version:	1.0
Description: Concept of associative array and queue data type 
***************************************************************************/
module data_assign9 (); // module name and file name same 
  //ADD_CODE: Declare an empty function 
  //ADD_CODE: Declare arrays A and B and size as 10 
  //ADD_CODE: Assign 10 random integers between 1 and 20 values to them.
  //ADD_CODE: Declare the third Array AB

  //ADD_CODE: Create a 3rd array AB by comparing the two elements of array A and B 
  //ADD_CODE: Copy all the unique elements of the arraysA and B to the array AB
  
  //Example: 
  //A = [1, 8, 5, 6, 7, 1, 5, 9, 17], 
  //B = [2, 3, 5, 11, 13, 19, 11, 8, 7, 11] then
  //AB = [1, 2, 3, 5, 6, 7, 8, 9, 11, 13, 17, 19]

module array_module;
  initial 
    begin
      repeat (10)
        begin
        //ADD_CODE: Call the function
        //ADD_CODE: Display the all three array elements
        end
    end
endmodule 
