/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	data_assign10.sv  
Date:   	21st May 2022
Version:	1.0
Description: Concept of splitting of dynamic array using inbuilt methods
***************************************************************************/
module data_assign10 (); 

  // Example: Split the dyn_arr_b[0]=ffffffff  to 
  // dyn_arr_a[0]=ff, dyn_arr_a[1]=ff , dyn_arr_a[2]=ff, dyn_arr_a[3]=ff.
  
  //Declare a packed array of size 32 bit named dyn_arr_b
  //Declare a multidimensional array dyn_arr_a as specified in the example 

  initial 
    begin
      //create and randomize the dyn_arr_b ;
      //create and assign size for the dyn_arr_a
      //Write the logic (loops) to split the dyn_arr_b and assign the values to dyn_arr_a
      //Display both the arrays 
    
  end
endmodule
