/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	data_assign7.sv  
Date:   	21st May 2022
Version:	1.0
Description: Concept of associative array and queue data type 
***************************************************************************/
module data_assign7;
  //ADD_CODE: Declare a queue with unbounded value off type bit[7:0]
  //ADD_CODE: Write a function to assign 15 random values to the queue
  //ADD_CODE: Display all the elements of the queue and size of the queue
  
  initial 
    begin
      //ADD_CODE:ADD a queue method to reverse the elements of the code
      //ADD_CODE: HINT Add loops
      //ADD_CODE: Display the reversed queue elements and size

      //ADD_CODE: write a logic to with out using queue methods to reverse the elements of the above queue
      //ADD_CODE: Display the elements. The queue elements matches with original value
      
    end
endmodule
