/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	data_assign4.sv  
Date:   	21st May 2022
Version:	1.0
Description: Concept of structure data type 
***************************************************************************/
//ADD_CODE: Declare the struct with name money
//ADD_CODE: Store coins as type int and rupees as real

module data_assign4;
 //ADD_CODE: To create the instance of the structure
  initial begin
    //ADD_CODE: to Assign directvalues to the structure variables
    //Display the values of the memebers
    
    //ADD_CODE: Assign values using the memebers name
    //ADD_CODE: Display the values 
    
    //ADD_CODE: Assig all elements of structure to zero
    //ADD_CODE: Diaplay the values 
  end
endmodule
