/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Priya Ananthakrishnan
Filename:	func_assign1.sv  
Date:   	6th June 2024
Version:	1.0
Description: Concept of various task methods in System Verilog 
***************************************************************************/
module func_assign1;
  
//ADD_CODE: Declare the three variables a,b and sum 
//ADD_CODE: Write two different function for addition of two numbers
//1. to return the value  using the return statement
//2. to return the value by function name sum 


initial
  begin
    //ADD_CODE: Call the function addition and pass the argument by value
    //Return the value of the function  by using a return statement 
    //ADD_CODE: Display the values of the result
    
    //ADD_CODE: Call the function addition and pass the argument by 
    //Return the value by assigning a value to the internal variable with the same name as the function
    //ADD_CODE: Display the values of the result
    

  end
endmodule

